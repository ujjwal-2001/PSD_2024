//====================================================//
// File Name    :   TOP.v
// Module Name  :   TOP
// Author       :   Ujjwal Chaudhary, M. Tech. ESE'25, IISc Bangalore.
// Course       :   E3 245 Processor System Design
// Assignment   :   2
// Topic        :   32-bit RISC-V Single-clcycle Processor
// ===================================================//

//--------------------------------------------DESCRIPTION---------------------------------------------//

//----------------------------------------------------------------------------------------------------//

module TOP(
    input wire clock,     // Clock
    input wire reset,     // Reset
    output wire [31:0] RF1// Register file
);

    CPU CPU_inst(
        .clock(clock),
        .reset(reset),
        .RF1(RF1)
    );

endmodule